package pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "../src/agent/transaction_in.sv"
  `include "../src/agent/transaction_out.sv"
  `include "../src/agent/sequence_in.sv"
  `include "../src/agent/driver.sv"
  `include "../src/agent/monitor.sv"
  `include "../src/agent/agent.sv"
  
  `include "../src/rb_agent/transaction_rb.sv"
  `include "../src/rb_agent/sequence_rb.sv"
  `include "../src/rb_agent/driver_rb.sv"
  `include "../src/rb_agent/monitor_rb.sv"
  `include "../src/rb_agent/agent_rb.sv"
  
  `include "refmod.sv"
  `include "coverage.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "simple_test.sv"
endpackage
